module instructionMemory(input logic [4:0] readAddress, output logic [15:0] readData, readData2);

logic [15:0] rom[31:0];  

always_comb  
      begin  
        rom[0] = 16'b001_0_0000_0000_0000;  
        rom[1] = 16'b001_0_0000_0001_0001;  
        rom[2] = 16'b001_1_0010_00000000;  
        rom[3] = 16'b001_1_0011_00000000;  
        rom[4] = 16'b001_1_0100_0000_0001;  
        rom[5] = 16'b101_01001_0010_0001;
        rom[6] = 16'b010_0_0011_0011_0000;  
        rom[7] = 16'b010_0_0010_0010_0100;  
        rom[8] = 16'b101_00101_0000_0000;  
        rom[9] = 16'b000_0_0000_0011_0011;  
        rom[10] = 16'b0001111111111111;  
        rom[11] = 16'b0000000000000000;  
        rom[12] = 16'b010_0_0011_00000001;  
        rom[13] = 16'b0000000000000000;  
        rom[14] = 16'b0000000000000000;  
        rom[15] = 16'b0000000000000000;
        rom[16] = 16'b1000000110000000;  
        rom[17] = 16'b0010110010110010;  
        rom[18] = 16'b1101110001100111;  
        rom[19] = 16'b1101110111011001;  
        rom[20] = 16'b1111110110110001;  
        rom[21] = 16'b1100000001111011; 
        rom[22] = 16'b0000000000000000;  
        rom[23] = 16'b0000000000000000;
        rom[24] = 16'b1000000110000000;  
        rom[25] = 16'b0010110010110010;  
        rom[26] = 16'b1101110001100111;  
        rom[27] = 16'b1101110111011001;  
        rom[28] = 16'b1111110110110001;  
        rom[29] = 16'b1100000001111011; 
        rom[30] = 16'b0000000000000000;  
        rom[31] = 16'b0000000000000000;
        

      end 
    assign readData = rom[readAddress];
    assign readData2 = rom[readAddress+1];
endmodule